module cam_mux_test();
	
	reg [1023:0] all_data_i;
	reg [4:0] index_i;
	logic [31:0] read_valid_i;
	logic read_valid_o;
	logic [31:0] data_o;
	

	cam_mux #(.DATA_WIDTH(32),.ADDR_WIDTH(5),.DEPTH(32)) my_mux (
		.all_data_i(all_data_i),
		.index_i(index_i),
		.read_valid_i,
		.read_valid_o,
		.data_o(data_o)
	);

	initial begin
		$vcdpluson;
		read_valid_i = 32'd0;
		$display("Checking initial read_valid: %b", read_valid_o);

		index_i = 5'b00000;
		read_valid_i[0] = 1;
		$display("setting read valid for first flip flop.");
		#5 $display("read valid: %b", read_valid_o);
		
		index_i = 5'b10000;
		read_valid_i[0] = 0;
		read_valid_i[31] = 1;
		$display("setting read valid for last flip flop");
		#5 $display("read valid: %b", read_valid_o);

		read_valid_i[31] = 0;
		$display("clearing all read valid inputs to see a zero output");
		#5 $display("read valid: %b", read_valid_o);

		// making input signal 0 at start
		all_data_i = 1024'h4958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584938502948371832;
		index_i = 5'd0;
		#5 $display( "for index 0, result is %h, expected 0x48371832\n", data_o );
		all_data_i = 1024'h4958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584938502948371832;
		index_i = 5'd1;
		#5 $display( "for index 1, result is %h, expected 0x49385029\n", data_o );

		all_data_i = 1024'h4958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584938502948371832;
		index_i = 5'd2;
		#5 $display( "for index 2, result is %h, expected 0x17384958\n", data_o );
		all_data_i = 1024'h4958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584938502948371832;
		index_i = 5'd3;
		#5 $display( "for index 3, result is %h, expected 0x49305948\n", data_o );

		all_data_i = 1024'h4958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584938502948371832;
		index_i = 5'd4;
		#5 $display( "for index 4, result is %h, expected 0x49584958\n", data_o );
		all_data_i = 1024'h4958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584958493059481738495849584930594817384958495849305948173849584938502948371832;
		index_i = 5'd5;
		#5 $display( "for index 5, result is %h, expected 0x59481738\n", data_o );

	end

endmodule
